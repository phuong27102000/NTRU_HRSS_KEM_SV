module poly_test;
	parameter NUM_WIDTH_LENGTH_H=13;
	parameter NUM_WIDTH_LENGTH_R=2;
	parameter NUM_N=701;
	logic en;
	logic clk;
	logic [NUM_N*NUM_WIDTH_LENGTH_R-1:0]rin;
	logic [NUM_N*NUM_WIDTH_LENGTH_H-1:0]h;
	logic  [NUM_N*NUM_WIDTH_LENGTH_H-1:0]e;
	always begin
	clk=0;
	forever #20 clk=~clk;
	end
	initial begin

	en=1; rin=1402'd5741759847443523486915852740064336562367643230359378364070146297719661374989682971036864603408974334467505944949513190067471921428371033585051426379762408058199425673207531662411762503887349139456528297338700945905778556785869616719856381777515319629774895725691427009624386999801210216166522177507739854634912563317408249998208898583346827077201057314384101813413754822716083231484489878782375027287512936581840526662659; 
	h=9113'd14601420238058491397818467492538628636664570603192285008487023978165991533410348260634596869542563664175958562439450911670204811404773878754547475112482130424019971961969266313811166599258650649548787800144670807924936876156173023062548573566754325375982820947594898790316284290847375945131608690212060099607940339130596682850209774524389931750626773103982426345213176377318918684030478812239272034919013503730272524273674467693315531084711815830918909826276840284267957936357812760278319727486532739854449436728934605462960336511781472235966223151434783720865140031360392517962845283467211966454105642953883578343030219746931303841456542404426041977896763832035888744617316188572809350370164469759666959339975304024421896349430103113820979486559390413542006692557713498424071676100192439275891672300947352791873030485785648205967041945451802918154383202132811960667131307305818008595537955049399923191374088269517310558175275352821758230286733503079820653659940433008983313197589427596055357680054211837123372092708482043669188318442186012871756901864789744038559268640097373827800791902212806661491659081671033468852508613963677795012857540241332925331802779884767501336089928525254092643894801185595362401792523108878921188228942896477187928752608962466070830344100321410600790058249000237445078406001103445561350824782155170235128576113807164374716244981889829007081834456523995945052498397837364967138683298638257408574378039515378591092466283136604260735407756069113690272487761326988818282786523393685471938900090421066638285736896529552785470126362196089829689497539896506824308095713591737826735206592691878157876669402130666421366777205860790554573060857926028131982286265076872092213912777553234856956800138505274318630758112773095370751099469729515596418586009012469527430076178187087904620183542889375880544915907640557976876917458969310418188783843228249246318476581969262750658845990494977072652026624714861449634287502186899373562242104033630559193443421201266589906491983091211723085335079099883322925748288260577943477918381800018387184427764875319201342473235989432084405680437842282918312009276173737653951564335274969343795261158438269547254385740008142656491630497005621973592963542289228697832137777679551029704746029696141846344464949210304636141490648172713857907484558401607585701709516311012780148881159272075245747530729334045421828617677612855181022022182633708397458380285381558856020875577877749201090505425845818141495186977167533101207136264641139396508250287101816012704123406898897191247850488298437542141325126479993167547296890210463405664737760960389756583089350806404449822265441147530946965196164707654000499732051007340967570737715081982425947045931065434970669746597539418592428682886208656392777553846;
	//ket qua e=9113'd4312971603255676855114546619287656850335658274688583909803132429324845082916952374051967601880107339620229453889904697707085107077642206380802103396710853745174002373374767578270260306340994624513323292666246363189792952521201547821516712191861535232587431521102866163911545564428833388979124402120924969654422235297863820832849738083370097175185858729301861181546346683850723180457495784677475223430878102360720805864184693087407803480980970614297487523222995653993982775707992498971678801215392509411093482758469294683812720663135369567337819979481909526350080048440399426039987204566769579542034409624226058635882194889968896236966523589116695007837643497390237581104201695127800382586803108388501626922693905068542220564819620253407034374657463982680761518247177594626080558848775649560802747166556780554913196793287916522043641976474298124636244844918242880236897186997867505859139792067831020132417455472200188301377843899967223499685012947366193911376200802730677498114585088755431386403139853354278151081307265232180999625615374118877993695102032898073031488315571112398649769082080573568166555372514979444854436014223287223788908769457861902916380894322358146535396166902742498662858437685247791134039777907165317404329879554248703586587602200687614696170316325641771760593947139705662408903220964959465419276820127658630600244410620145992290628657172337484875779849754876116203864877472989804824275116655934075429699778121583739929767429004941709681343758691079440977063191059494299470104023504719157267746924443296978804569968363292009117014732903626075386142135911648627721316624800294191372763319451004872381612477925910949576049562167679385167681735144716305166334579452962249663711096199215262802625757576932871805788448956724749008390752005142051228430042363704831711950431180747149672421776639621841135527717753075013617879078587652831133441833441410174177431817659949969425061840302862261722277364876399595616523227638198810622080800657205007278159396431680740734253954324197819395560838143551726938322650638640731494608831060400810566781054528187755744142742679517030025557597285854693791585835470946478712620238717818205466993243058071246769949635209946099614451796655275396421107110195050294002799511723282997985594073307348275169366315623818474385100898546908283829527503170041997142757413380994630581683974353478551465106457596404703073592534596347873902690097114028978591217168571957379875467575059156017837709986291365986227874504016495690078137731602990413299924066250058244852849506919994354516641324524952128183239884601089164921611409806764368269641643855545139392074986794879265308661183708385670926560999355811341458142912368602414564870157922384398386119412725053124113470737700385670446754602022509229704213678s
	#30
	en=0;
	
	end
	polynomialmultiplication entity_0 (.clk(clk),.en(en),.rin(rin),.h(h),.e(e));
endmodule
