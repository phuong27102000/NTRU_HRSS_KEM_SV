module pack_Rq0_test;
	logic [9113:1]c;
	logic [9104:1]cnew;
	initial begin
	$monitor("c=%d                    cnew=%d                  ",c,cnew);
	c=9113'd13489446077744938222685651298719558073554355724181941307530511843429337676002508975066364227363667444300691575548118192645784041629033652457597971663340160872632967012292707415005178854021391368721894941015417252048937644949012095880173256968582551122919247023759372902750551686636544614112780117075839526229524179478489932513616090989041728302545008507653288153259067339330109693689437515503077179769582257626668636335525320682164004583682594528891715139523871060745540441892176538907268061509234249852954038961189084231902090447249910552360494625216721691512873257391964788958087528697562299888575437762901669368283258326070559037986682414338264286382528843166596403119796931307490966609126013766036650383203085334495217280881065226216249392893251204827723108157127979145682947859931784014526012761569961547870801692654227758300252579581510218202056831600880524797746809734384383624341792753248290765924677215168916133915827774336605046154038045191445765317014706853623700857121142018822729279439992074520796502352535581305586780677370479702011157017229388849320809910382076930539189888208095294264656418632921625332895387851551516309152989533321397269396648409675725573334296190785520396297018425176355681476404932703575797328424487220308389187638382824400345985937129857873630888233970400097275213477505760683583989752659674668877074765627626345067378274558450172410600754590105766180511185171592640588602813380842475438449060145487620854111210629156743136986312727335938013437309112047642974333667059641607528389625625424674861434012336019710529888977858832675789963671215500129069596791128120703716155440347039378138511395008066816746094712678670349502811349504209662343729964352835287328548846238503174884686918606248900052414070164395488190277165886935444151458561308156823784576221308367944647839704295202347301336411327411441562575221510560685393630006491170211300834426659298903134387926023864039549549248897085770732548672565329255293999715102276231392011573476266294425268434602195362309470047859096784306133354995701969932300026251063335430811108716358021541934665657586683449751295177819212102952866856282656803566006988828575925609064331760389779638776985080710077780806000182447934413341681528864800946236068980319772972493264713969822822538348034192824707880440041558897497711746505909229512198314267598449265258740110116569950084825516901266802246057678629097278361275379730238834045083497846656942837833570955900617280546215891734549588975157334594005215055675724693887054785188274681817139325405410707337300069187767533108807081806451007723318915224622459071735863444755945691343924171522456391321475474977705376794962679844310593207546598255050927361774941202934498706395600814360987325119489022257640947906788614995435616;
	//cnew=9113'd28381927568259374097798126705792370461034790296954733358976679972277706666883039930893032764508806003983243355544536131532768941232249590828586528732522158024268910940221251810114343442176312020859551129870445473636720797667179381507145577967952050640473031323333007213924305189106650430831944153562376025451507228437256557734824510753916731441808153961743965896997589562365443940233431285965989357380398241059915580190682651932894944988504382804618130515034924595336861994774552728498780536003204937462532398191747858336698826280203276050961868426413278048593620338439286542896447065841356084213552094247288294396109378661255184957476738345586823374356537969678431744032484036762951405315414302110692341772742850898998108964497396826402381754806270769530130435469271199919930523191442188591169282068225916844217505063775060860078127157590704618724503764805082228048357872909165956656467462743964677852568302178731369009799934034442216126433903027124061036179674220364026153607057468235325054115698237504211568377770356954221247173787088302091675433556417605487536123739842880122557787726380688757141228184531313639652850390528318933590130689966548824451025848770020715907179138967489259558766129344625371138074109239657366079316726417845838690114096354404226430232137431929835530901468861846690871680301836093377094354120277798695966160892348431189732295018413228682784978972953906151000175124552725424445965483594074246293749310839992248950266602973194963323980199186849879212396785490532070217837050859548666357597476016699817927544353867030322336706472108501648737002724958086014895034169515799381758986064962104077305029450688003311302400046100559568967097253654695271373434235476123613410526429833391126030551175198817555674263602439665627177844726891936909769691708643763631377876296170188204422421757130984200850435288793089644187053709669195732329628026070011180450055063198084903608379247422764679353284581029427929908273696133754128494501852501838894196006786442011539132530633051292633418232511796709128039975125553983945613099621349673589389567246817396159954942986810318581907758710212513072670663082754836145830899759760849701386357487477668883467681663921029755723216340878728171356304463488149217519908705082551031004271417960089951826042393667532147865371343247739748233775896493254620257542134558757641889743452837688037754262226134919181770592566614506511844862956965778397351677751822613457019711543051611784503247254969686211228848801301123482579664763294560232093519653050325826954162070670499632340027151136754612806055638528884503740298671107880328831908846315439258795260296635778718782798224911323483351999039496187765843349598488827353655777107090475405789621902806002194420474703009116859771821946278236819818246;
	#20
	c=9113'd5290642969891323020368168308931744928767849464102667205252884145212213642742017652342229265455562741034338132746149774905188159073865487643726022352599310487651268511224797661470452176351350323109735533356891631287875816885763828985151082101651807701597604789196338864114659187663265400807643310431276633959454059622365366917690463436595534233412994913118386606824387201837358524648306660416553918544883695677245260513303541228450831492800136164253759580243265744827125109802956972121757416435954502389582231294253182730825939400419280311088323903050457789809427962664750432231426190407109532018843792253251755539108231365041550552668709964070856500011426676285849082041909808364749664068923291327651607411037235507074970164432714081111407744626999088991587153964088131966073263757745838647539739470479545264649392272726312845712680342556297386227747617910423104456932927223579349841049364946698293297099361813583536405001414431483380121945278150162213988196721304324099538301483072316330970421530100966619146550607658127990812369782170813853938389921263798309868321910745803394227050922528246403148063167604486176076093471102904386634171519693484455284620032981024635983770003070146383504390864561703153671624954749697445386089797198348581398130173529607571949361639554724535044958785957784045410085589603344328219605573739162669180499768368467068289627626663562496915586067884333897969256232301283783312699004132428689824858123878761491976760136959033870780761340467900634748468865084455321268946815447580535368395953340970066107982921712798990152901081918439667815975677614318548239145235338791784224687829373619532120934821030608776065288620851326785629499497263879275673696356328154816234235223299967779299881189398563461932506024924991822519368252357877810124015440497489639235232791688400832331245711572986570595148125225225882626579984763666748006963733768660869794619509700054180663271617083315677790288495109826237804095412953353821329702104736378051176634365981715960281463691281013517195055966679609635441265278377224121259363649164441054814495316453906766361694131466874588303841862246209004905415214662313180421452316945317437235775067176171554664185754137219866888848561203183201252569110595022214421876408833634115288009565175145645818358929663633355007998251381149782406327132910823327733570272272623202063033463647697241452160159167730982431595925066572223580145686732072602882260011928510019153003345213919195406404642265017985286417664198332654538605497707302631750075982338399815730833046629267417338335628658850174414461975930827309897682213259743702927216531298689246910632252881046059191854313786314966195840198831620237161816668208814500715312272100257712691464789980631503142442686326053910855273133174230759904755134;
	//cnew=9113'd2436101846895963985452053333992090793416853956113180144522022563356071569766776799312847827001590797383027000072797721592169685283547058101622699405221107424326999626022658747146878802825474171037202754579897912160489223199947717303420932005135456524232687200764763485149085965857765111181239415719149892201857470353411124285856672706947365500294662398957456341588444276713561577547788601241311051158675936899202204476751193628756092180760335847551610088188492610606624058356734297154139115272854264979976925022553423630072441270085767047256063287743420779112125135959915835114920102891116432665517207235331695060032536713602933319105263530683942708369020275267035320312408511640603269067485053501431793519445636799970592318565710089273601572065479563201288936695005237901208342318775756494390135065936120426982026958265516336331251780116301112522175366347227432125790277838442789182880979876587537331545345151792318934192726035532764082989546000389906943067896125010635349627963321418034818623802067742248914194630720972831863449077042495857349300680810099568888942899624568819317139259881905195923294652045462042395779682731877351895552415114461744184520017256594739699071012324445377624127438881853037214271111809911028423070584722315088234441597063354355557839440980852946508056865057849017251406423615938925692203062082666291825722540816069354947518054096447179904732801630377067050883187697295674241777925974652534196161164308740152774614009957833826900838701394967443020992628859656540135731271983504471025862507226942598694237633967819501486708881928857866054953875914458326977947993349098947933008755765109291146136077497200368200555070558729953237504107246030948094736932939922429613351466020684122798896258794326934527453512699198285848928384515690737917769646178708406960252727585054464370991506044466157662255778681385429292073217838878038139755750350540336573554364561177853038273180691864469526699123736844541401459620758946543670849683800611150761857412218072717453104772160307704065683709919265956262355750543543838058285200722335456615377016687356215464895982463237482239933520683779253921782647958604829646264035928793241530456705351125780460671663875303378027165576738347158862369189296374791360089413273966393199652230912664453769930349214198480972765702769083434027533259244314353554602180746569043245186968344994713815786584867216918669828784063464793328508439532952699108782010513582077449286730427395977700419090697326792114756869188101718423689318931985381175078841624815905727338040099660401860950406154104409813824637680034969657780646060612376688906598017975302494273798646051691013085237299232164796865873625918936501634494397370031786813953464581042761006361443494317165002249793049954311510606244033098792317;
	#20
	c=9113'd1560764698316765654979052512093627629039658012855778129922451709919379442395766266118453590649713126949448472773059901039667543946273808171737053670133270249205167143802402672942223005188409040514790859303876175093425379887353755640278071637412607039938984773204938900216666872593702891474165422963654520333592822391855921519074307423006603008374628861168378462324741576096900984344008576449076555491922589622036786649238638394276110737896551162339576782854235257184448486987412114584664825863403131614593268237212533873201247200857786116085944808867245711924292953225690763451208995233214014710397758939917697171929405651881956612262582986605402063718935293114887161366332487451078362154117894876162540321689736828163217786589064625055302153618812044049235657451822660275401635482280004409168107963033702183446771709311799725676726265320983163290372416281631988533390251289835278527451598901155201362196556554172281391480762474493655693140200160121948655964052053912288914999855534395663114102449935232775515272190466321027659730643977295702557620582055827083703094645242569575463468078920643296406447522019507398532108475868777665884919805464128452173920949942012502523625134102081102229266656828632674435446465917808652747162448760043010011436115250643957117260229693799736595861532893156085619473832740273449329405468988148360160865135409341343822904449181686835899641787020873597678688174226104002903177498274625470297612074894562345459095881772024595268290174073909246246943180105881903303045320959048337006490582675942621180557888240032711089862362552442305092710530813954996254183322646491401939670164089722045087525903668872801685822171806775700178526757934375333928762787506115382230265886009741449767172530057477136460542940134599359866917832792372040407601896993889224302631513499695758414614661507082623591847854942603697336301650245581563004021874513836303160605679988805435525195384460875001493098397579737199460456294174050472310802206191371734441576329195669024543100881813355551177189041188585752201242041270970358411660477207460756054200419636902572848206630356828846730926699284817579694678245674880018754365444904015367337427225026623120067336552083872488539460671287539714691183963561751259295020490145009929600291121220011681171887139009082453128831902871558828687075986868072870234770706857080476832015852472785271741544610389130279839031651532390568991442853492566132284800385508306169888452081591438432137772913746964112117727446438724310125305831992421350785572599618104985379969870283142020801495636699357279300018388485778590652805573880867469675906044492670315046107387225589986730298356079356825518982481073984542679734497922706853194784937363810470199341614211465125892616401751004183224121279288484932400508505;
	//cnew=9113'd4814327617422915703962863138549501641740263390330760191440714610765902995856376431023160729442265634362101261024604278331292142563238270041854625179799259784309954410032224534950934858041870877163270076088013751988119750845636761355008125583822605148104045178883868575401897468381884623944025409014538076580860133450848437160485718442719956827718924045872001575917202932194421618570417585671473705151238626779192317909165578513783039659105047194778835567456678526532740292071015169114398174629798230632376950206935179417448676112125597346938323083260617578904790109979667303394837108644277860001238303604137596197974423489666699068529557580167592378855556193451878263916264875071530214607077962326011616670653752728396582287213561968544640367278127583515317638076794734799457061770305498487598149804075134329020148829399713613108459858796068164814253900369226937123040401901677015037550910372776783353788068151895976027111678059947506849236387504844004230425587708363133353766007502420875131773539104600455281950418920953388571925488439872216235565376997799310252115039836238334228501905741299091131778687931360012811925567215024110110585632113319557523564989210776171208061234289437981121159700183415863941891993991476830600164939957779016394945176887230946473570671269291022907826937936359995466877412732111650970593092796916297222165962063828064994035931390322849340665308168459528783819090592121519645060986791195721034051453230743718126378718947978488324009076549052386272639275979662350054222489441607464715023920884754939602372278063746777952154021215909050458134972725003819067885417840297630595193559922345480201692095317234101922878259957406715804454996240771191573119122204183294648313482217739484712049121081392319145515639698937521585689061656031160560939500632900102933238554338924614060203854906592606481449652041105312502602005514598282378383971009581129144464604660622505164362790563328645399374399592265792761128115973525523159680677771192017714247955632424915140539835705277121407113699671264577908012051986066968828866926180775413399302715382579541947496013778601430621428785259528766125133808513011216843028822799537097036745241231750493781683455391514398418298890517658148350502294694318940205960236121926220846275591727805715967409080766832270799482295481373827839249439500758786685948952813715246790633829807760574521182536986525092566627515013311676583554126295795654155269996644642928450075800878822440197665215120963624728794438826260637112517480458344006084716848659662607605529245252493873286384645387294267016705590630333410441056759209861970254731225196131280347107790526755314810347162225412351123816158486496554150578050894717589831498105538839920701849786928177108323678067005256015769450745482931660552090
	#20
	c=9113'd11248618102391018207654938740692297168346188488546597299041082818469127219540670977999742510715693437026927782595315253579500325083856672779240653511467022801657026035388554451083415745968553483917788045918896698713559379278017115700050659924374657926412179118606958238657233533748922526480633876408614938821702501882609894416802314533241671463986660978606090406605701596068964996609989242828495491199935364375358366846857944610300018113351200146494367434219850050657642554528303555527752515516341173407568887614786008139443352519033816783635537646488024022863773197093743358777499906658714306438454319715350924152594940472980022577716097466156970889887236151995260661807582687875674560164082340109791032652996778589598124908847850098685026093516179325940400638386441392021817896752380309557057215698959173589747517765384655760233031284802673260775013100103671889691513616123984155589330325834597628696907157443041097447287308956170767581677643883013831982482925100434975056546210195435869725103357007494672811982397106719062318165361359419125806138168620865170749376206462016968608044166001149888932157765410176392556458351898809226005704801246768899761909646224143062829497707107334499496699839541601475627449465740025972766271612839436661467020666517015316899836018027999102365654467792055000379829739023369048423311501390806010046249391713577714862353639580486420690010995450695004938169304137767344448856914736068800637942605055334603209737697375545899418344987052707954162441766186048280435767001496639513230721357642374060440452039176027473340767407216504395068427480734178638138074826674141897173133078766137499458354536929754852363711530488779185007968558721316700092427147315734300956628898393170469916399282573468155260315827132562834232527108540378757166304182405829172500453559935631674533109977037297852273896311343560104206561297216448598337731276678288180251363938520951943307247068399365689177200463370887167035631046807649545231089657085025601746550493298844853529250720305408309359587555214679790605176809468640945785433182830978852342552581888032128556681200168639795288094263847778656711541266187674305397978473810712797938079365785784909585874653125682987864579985064853912780667941329293245233939402099207504430627492143174534345193512543048554091172516786320202370350842662635011361187708472935487737760997790022209267816504766985582281770897990050366362083348403918949765033961277135068736217727709984037626969192490876081475452513168822104787308985450244185556341436960240433699761842460771749141964903665462888829397462588785511118236154309698842332273739060758274303575474303771086964816856334769701892466607864312168551673414292749039822831810023625545903764204404957851211334054701637991208031265914449610954444772;
	//cnew=9113'd26084177933187962087152022902130338511500220000056897387116757197848621306000013162461018010427568457435951248353463838815814257870323548531215713281258179429036771497144497106490048986370563967191615411805930351207143342685509968498248345851202748506716421494991577399382149016594811830755733671863936813304603990735743560718804788845773057530328390451573683172023038373257411800887817551311942151411979238020951652376389022438841119385409378148516943085475711806524621075734647350890465854109140735304151960345594790227959211729785068277803278869016351823489675098883394625410073479728885661826732581312550281011147643890215186551004422161334544733639137678209028368165736220397508041117461787534695377769745408652465634509853783616977952900183346812524699748505191901328253196925990655661366701167751666223101578981003905928842810836883911306748566043257636989028474916799515578861284314009565793381959447571535790427241125488963061930582641757909914970057550310618006434180635507667281648696162830975043408572237271429938514057898505730729401086251116737969151333417688047500536943048322046561479863200787349248213116431345111872898091099899979266853883383345481671905522163304551221313946285071403292675548738780200744203721747718229356393279537662138042170041831486409556965828639101263438203184209079724846175934466599894008916819825103352522077760587198403097935321668729903699718094456063389963124443669734813125621043794594050772920913611880303679626100405415657770923608468972970363996943526970564535977990623364366350017687241712490719886029269050160600835755214375272673777083062877176177884857864304144995160160542465214054052553799709391193476437980914430338846710588210509942660075393205657880784605415003995032208910959099660747576425790329184354139912197397290119930703189471275717846117928180238311038225752542405679120427200015336671871326030090887113533245529466171895350500505552124925943598622619236639515548868058272653744765965523833917660981289500665718344072919610088477742963452547792500077264752403611817435197547743002493983979367835910030213751898608225337451537796702347676025673278345958047807704722450112784025997880101011317671741568613002201342264069831997087239168879660708508731611730721099686125088539766719639362566106268742994988190604480120374662172394800407492700980242274846035790907346905827639273232813664313698714617938090285830338006222819265405857015909037339738967654939757888774555170752183026344957894740020742048437100057898247672009718930132303383752394112927811897827735699994362429670648561314201055821798052098576703478760852464295273499185338041479238785561123864307327652623732496062320749848202598259598407787134358842343467089975344077926540558301823587762522633262812273780191271;
	#20
	c=9113'd8655237013337022778752977145459788870580288785088551232369038259706813724709740935887898167551095190020688432082137624898861511743785396004793645465487219639086999518420748425770541504357479761455348642927973811988296402195433325292326623048725676122618885489005262933020236541754071523500313641106100529610885456117347959096846392419509696249464182531526344883240941358318367152370565956290998250340116196848584822727915172456818161206914277800502366375124144713687004618911840426985756176383589987145681476883200710406832724964631284875725306352956465488661129606840455892895572274632837221243193290327536075812466809557066663790904333784284238966296553035651044915259665574370781530713847628028944849229652471454241115649596568553546793749570693327834938845008726787798747194786418720438101501025911845032883582208228756245208735260989796859454735297248131769502307364719288407104190766671345818306581400352450244425570828931188442687091441938099627378929621906823931115911029050638061746306413754198420651088251671488074402012874071585069393222083560005314835281688561900189983957539410700451534207168847813024358074225486292042008354296381780857233398198471545081995882029938047957593083538781727000196747112768816283569659054916907222746389566823953717351978310067495927390143864669065577959713756444476854577115526109182298211819840728510968460481991545915664929875194674578770540104882881229039268978860232059287102182669197584867802334442359019351167945233162446817524385458954098661745192684628678025978168725119492201556791759671609965371488842683627662675120202984899393821749980553824331963391196237805944355846234247618464394689240433679434115470255779746006465670091254674060273645387708581122277700411442510727772308419593195836886500799991679361410215301770201819894212234808670331645500098418929102071986453193369045140875911395709055649735928482266739107863265985155254653349475667982408570578082519084092162101808186097979022501327093236099570948891245372307431805356209959830974702001179666214908433294913365059553014125922958083728044945113487039385759951942524419356901391855340259817881242201194278224410935707763232631767478569534970270740445675256620182140185127875347410936026467889746863165119948498640689659709832718426922732204565232869118294278555316242085520940085745273850818948708280071379491104167499491868617869338455435521382441406558236276759942626055974724748503014922389962729846550409941280418963369124749830353176198248526585629167544940452887742212568696412632227816545664958302023132744848209131049835208776883502869568552303943404267356163338864049636313876068299112630191053252297180854244337610395970422469813234384443576997124910920613014488305767576000981521569927259100265310323487074035343613;
	//cnew=9113'd18993133869169923031181808338158726781666209838948360272678359605369005728807468223536476037573790702171818004076279906778816277534492100761865559008658608394096074465536206566044588317960115905891499437085114403829549243695511612942645306320738098057838057123079047471055235498521907681893666006560454021731349546103220602143376814769629654347201573255228056465769182753445130244250750554682038651187282229377806376230723975273588873386130212326084925760043804918697008655985523155201270653465110681780940273592709131821444543212992179276628466450372559993460914126258870564907695859427627947107831427456713028846055158203662784153639479219504920438665237441978819556039861041145434451553391305150447944933067310366955174144002650685382607728438324455877940220415245101503580813745560691290706224719877419491011399124635131111484808446164224988342862332555419262315944885112370549973051525403321291732561903050915641754756611977162850781096229112109138047136411170049434105231219085410113564971321785805588705925517555593003701508783441402497957357695782992725767213997806314068468987663158443097493985147876785341603136335023087575203424755687022169225795722527254645778927997558909348017814876660235724938137717065598498983710685874619399992537507516655544085986803509841639669002830590381468365588743948309779371443716553410896571533337339286394860743743746897907255342201784783635493766493990324397965189942079883518798053729078694290792765557509437615061828441586978944795624520963906258775258986864288502579075452511936741211583567485118832039573405837000658984631212940498552736565263688381832612296583655758024101365008442910561257413623260620883105048900948436249283280068724599180179589161797203262211620173955358781100944098766374721548159559726191798102298779393374922003328776323321648656805937589157539744378153225444021170487060318694831424616065301893591518553799359402797046666165384331714258884444619889401355152632584062905198630380292334726387460978180794964990995011749759915896937878464003033242078023648590885371767504093877059269969638617823475026306410021105412475952283605761021637208182478600958017002738630090477235124749485444624594405962718833441298163060862633292158547256316708922369762878007426830389347761431983542805391281566299936535343958995107249361942401315667886418752609374216164019432715579863141812929153327728825294485212918288142214973676963955910449968303688834004266296101198069922285787344204768430154051605044247172185253254229873653788668248535691362519276733624100354812210742604210290160646389027843374637956480530038665908095819668728165136341963766964601879097392269091901063743705340046716154778174007960903313648366346921170633984503126030746661933561763604990290963595634038617933247;
	end
	pack_Rq0 entity_0 (.c(c),.cnew(cnew));
endmodule
