module poly_test;
	parameter NUM_WIDTH_LENGTH_H=13;
	parameter NUM_N=701;
	logic en2;
	logic [NUM_N*NUM_WIDTH_LENGTH_H:1] t;
	logic en;
	logic clk;
	logic [NUM_WIDTH_LENGTH_H:1] c;
	logic [(NUM_N-1)*NUM_WIDTH_LENGTH_H-1:0]h;
	logic [NUM_N*NUM_WIDTH_LENGTH_H-1:0]e,e_next;
	logic [NUM_N*NUM_WIDTH_LENGTH_H-14:0]e_1;
	always begin
	clk=0;
	forever #20 clk=~clk;
	end
	initial begin

	en2=1; t=9113'd10668850038505307097012790561037827119524514281342774960634266848833313619791030671956200199402391694917975749057204781133836074973848489132638030198417020581517831888731342067666818407872514608848635789338818072883898889089437301020586372186657679752135540593613733088202086967223629894406833739848393308273452439708582889166479539023669225541403711578767836354218566469163041501032132807358039801618741453028895105755783902149729565133176452930763178175771506831910030911098351473353010955243652003822714912440430143479466119660300353753157323330414019834289132266520463811575841383698480861758950620197111648276629905445944958175501406496213431059800320335867980407958215770133529406254524541829325918590557254715090142963645527005271600570025195151009549035921174142689471674717829228658590850735272772124931979721769915581853347278556990796147058866846968114665752085199715850985382783384792578244032207013285373470382701231204304205539159260951273361594261798978421814098490124437071575374945946026903984343609442779998624784191085239927770423325343550108582586619092971701962568735531960117167884197716288548630391337073067491180442650168686217164725371512472605458664702271124883970790430551692692869882326171860315854561847453372242364502003483994058603858984588155465820559613696384496168479791907167268891353598280457523261058677616081390189606794465403310854142492169221669410645000636450318495380565712207782326450007484006019721409941583033414621875557034020766198483717273876584822205027854867533463580321338209335590843503697578105682064851010942401986251117299614075542970004651815361075719143082612190133686649031838318469882707788340129303450722624472325653313378085108301778104290184961166807445341281563306599218726218186881245973100357319037433510088397758109901612284965834684233852659215775964692102709965409582000535198761373114364581300862519798681056722881220180830631362666360871767536125931171333555289383748598314046820204027890030057154721809437702437209331624769376167055349374354188941043402850906463374319024640123933274192606337537272255929286341802977779902228564565887797691554584590405931026616466731241168365009403438443904307594792078793898808176741648894522653816742127452222074256334694065864441863036189425411463736436610597086491686674858781897921690576362242540713461695824636224196357789623363528836447836469817070784490473649318085649634475277082094181312659501382785217108784094416453556821464316833029916258608634505089716417032865962373548586432456563302853879787841460393640557132074367941851118982855786229634722825250074744008419649151809758035417131221783825851580896329339173386080980803351480082243633573226033805222888556920072291730281231709210185812557434186524312354191396224396152199; 
	h=9100'd1756494577084631577829860676438761377886098958386121207834194523547318494470442222569338671608406564101672187562534213742683007210045223114593127368363705628810230801766423146161621677144508392854533013515037868897256567202824046434494135631728364919700389750662039858725710833605071658465039758456335368674211846777297623411721017769306455549645960736674060444477911064760489048007051454188658247493053397715979158715727498525162947745122467932141692819662795134462960297706138917068177231122818361224224157079486969819992404557779222716497594039067742678434718091178543589841994283167459048429544196249808817678372729632123316816676861153966189072789900510435396499766625842046478534411981931092403378359497820001153774023520383232514732977816778893831277059993201300139465424611706383360723969745163167603702492557048496248713856541330004153301079453047754693941102224152098833381682977537362187604032438124433369113820810368752365183635017866236737691391883860548909746386936463789057294702334608514234188559267001554133797208922076447688894883024961465603671761348006370248538904381669712930973009285488908441365242552059805597950948595029212099246935523490227698108960156249992945942106663606736604839448395270571724215034845361221081978317583770852479209361113736845151548698759205344573913042013424720245322474288242957324055485416618720715337482159070308929465588547146504075031775989205536733702344297631583421118788227306421902233899780319758971894170135778069127695484747579574114863499589325830790165131421719567608668051237636128512477732831616849631570783933153109015689007844037803409330317455334832206216271640081182471904037732949131852368587644171686465680981265772305008476925224489158048544269426104877907571067683344738750143993138249219156490501963875302237455118246402388630285973920252863882546317020529034773783281196386122559373248641896757106512458997690667159747135915635493981827193448743589416519477920192444497101520812079101795599783800234949624139964454046663959446772782109983160135331246765511660100743787420326407296346861183625055477848658063993237583762228710459050652621260172137782463631701042609033127274890921353228566110034287615549725174759243212703906735777948153995845627369268342135513936684309192136095057440520210747530719910650763246581735373255301664370728467812797878654609331565207051073453167731267029811211075670003356181055680722076237961343516769493653041117307719962816166633213139887932741513836563089161138017614960860109764601455656226591617056670802896253001794082913827921359018337642608176248250371614816564716314717570883294356069417172957750255914520886657603451184134916376357504158580684312557419398340808163962292735336504868235289029766327454779455927058315999626983044;
	en=1;
	//ket qua e=9113'd4312971603255676855114546619287656850335658274688583909803132429324845082916952374051967601880107339620229453889904697707085107077642206380802103396710853745174002373374767578270260306340994624513323292666246363189792952521201547821516712191861535232587431521102866163911545564428833388979124402120924969654422235297863820832849738083370097175185858729301861181546346683850723180457495784677475223430878102360720805864184693087407803480980970614297487523222995653993982775707992498971678801215392509411093482758469294683812720663135369567337819979481909526350080048440399426039987204566769579542034409624226058635882194889968896236966523589116695007837643497390237581104201695127800382586803108388501626922693905068542220564819620253407034374657463982680761518247177594626080558848775649560802747166556780554913196793287916522043641976474298124636244844918242880236897186997867505859139792067831020132417455472200188301377843899967223499685012947366193911376200802730677498114585088755431386403139853354278151081307265232180999625615374118877993695102032898073031488315571112398649769082080573568166555372514979444854436014223287223788908769457861902916380894322358146535396166902742498662858437685247791134039777907165317404329879554248703586587602200687614696170316325641771760593947139705662408903220964959465419276820127658630600244410620145992290628657172337484875779849754876116203864877472989804824275116655934075429699778121583739929767429004941709681343758691079440977063191059494299470104023504719157267746924443296978804569968363292009117014732903626075386142135911648627721316624800294191372763319451004872381612477925910949576049562167679385167681735144716305166334579452962249663711096199215262802625757576932871805788448956724749008390752005142051228430042363704831711950431180747149672421776639621841135527717753075013617879078587652831133441833441410174177431817659949969425061840302862261722277364876399595616523227638198810622080800657205007278159396431680740734253954324197819395560838143551726938322650638640731494608831060400810566781054528187755744142742679517030025557597285854693791585835470946478712620238717818205466993243058071246769949635209946099614451796655275396421107110195050294002799511723282997985594073307348275169366315623818474385100898546908283829527503170041997142757413380994630581683974353478551465106457596404703073592534596347873902690097114028978591217168571957379875467575059156017837709986291365986227874504016495690078137731602990413299924066250058244852849506919994354516641324524952128183239884601089164921611409806764368269641643855545139392074986794879265308661183708385670926560999355811341458142912368602414564870157922384398386119412725053124113470737700385670446754602022509229704213678s
	#30
	
	en=0;
	en2=0;
	end
	poly_sq_gen entity_1(.clk(clk),.en(en2),.t(t),.c(c));
	polynomialmultiplication entity_0 (.clk(clk),.en(en),.c(c),.h(h),.e(e),.e_next(e_next),.e_1(e_1));
	
endmodule
