module decrypt_test;
parameter NUMS_OF_A_TER=700*2; parameter NUMS_OF_A_SQ=700*13;
logic clk;
logic en_lift,en_poly;
logic [NUMS_OF_A_TER:1] m;
logic [NUMS_OF_A_TER+2:1]rin;
logic [NUMS_OF_A_SQ+13:1] h;
logic [NUMS_OF_A_SQ+13:1] b;
logic [NUMS_OF_A_SQ+13:1] e,c1;
logic [NUMS_OF_A_SQ+4:1] c2;
decrypt decrypt (.clk(clk),.en_lift(en_lift),.en_poly(en_poly),.m(m),.rin(rin),.h(h),.b(b),.e(e),.c1(c1),.c2(c2));
always begin
	clk=0;
	forever #20 clk=~clk;
	end
initial begin
en_lift=1;en_poly=1;
m=1400'd5348781957263701820311526337382083045908442384806069698511068414607085671528498313075590681518625920548145312491763101886640487460530913203329294545438391458024591194778533438404073579896179565548831300796310152025777671122464183737290759870916276084770419529312040186625877526958233137686459731508531847755451630842122875146097408090672203665760256929123737251807199498668925417278898272143061939195014862493132476217281;
rin=1402'd27568469577021766233920522815002879918457521068659531775499976885059565502103555381036876842492302482817622763844710004235396140591661541388354285384273730715843215818953143746573375415655139551494058776278136806677644479142906824013960147259162763091738788329453876011631697817385613986969828394761388166237806417462150435534152383000897813588244069515639748258303725428021730129937179608664096395200540081656389086433029;
h=9113'd11112300006419830981102813097191485995506379688865442614624356227055610546520524785672439947716934624459785133041210671318087892890822053073932529621316943348912526012168593387321342165789861875874376641124486799825288786500498921033851213679085090760026730572598305796395107267722055128849138411566303072169657776711795613844884006799464955192779000671598643726987640177638148793783928135945138159062972144852374898766057911943875108552134253766915219923067812726328667967804076384200814356942361741647781888367026110858292028543205068139978837291894480157668982277130598489634174277942917964254423420123504129842243702560320150357821289376505840674829818375770922839049511322541463915488908322589015770307228136396010371699833369655863387850504958755168642148486678423152325029721553680821359261416268360538645911772139687585458315722933657681042818991911281188009442009447079020396593834802236399697776269233702342491646885593224042109234891799389198019778227709676498680015417048951668227430360037476048337025804726699952447404106911821730366735404507068719093848799980734927395291388778873195518844750899053882188017782607385311403411679721313596239790856446634736613391595628221029128318873307543864065087237585206154487279374472157034162845806618491739397706939830439072544329403231944113886635087670380784010882346871886861422311928065168718158939403379130250349697091521621900097243981215540884048745631929894124754907129112868649863122873064292839051832070632074771241927068899910194703684611053961550428955634064313422496097887719126067322676992319653846588722156613487516424733195342225898989137475349183534465532590676793177484395184582981878098916353074207625718034577755063765871081351096779283821827801869881825449199135739222849005789226733665881693208497268408857327898367950807720600059998706513921302428199352152533928346823465208699368963895158553003155977331328923619711642365588851968350504463590713246360253781896456339157650381425311258204202025922916262591771640046985260192992734477072381943311622204682105046022537531229038795513621002478242022273652712606093351222514198892182566163835646715711140853877610945986979719693308796044212417207012237270564528550977456268930764460711221957405986412705284974552439138325661749501145096243674921107804996240614200448739846843315313238563021147297225583755021067742774700541997350782345301788758145349916445122410963313129316474926293411636844922326905678687892234614549267478550487887882060860459345519684404131748844276306273351715720125722605521034214977701195638114595777662226565233745004469806110106353137524701163207575244874732835734905007404191765255176557732182760821773891068866191519176628175712613414311545779527349088190988151660521644557596148244500583200720;
#30
en_lift=0;en_poly=0;	
end
endmodule

//out=28401682154356084799928990976804705974021034820818725402481645416404887070725307966203097990604549226335438445452424100174030813061952362059461384063458225699344882349182005525386070333063560837483090027190077859604249976590484564564952856635551797213671895249691303268197690572193643656293455310292054739756055103602343378711810400105441232950792314977409813093910756193162225991764262358633172224377972487145818332219317468806407610401765775507447842592338040672328567981921094541519296368423915633072193149107407752475902042288123658630378627787444265939005696703780240385332995034730067621290994470046026437252251334411482310264402842811965169009380675830563125941414515203157784384066044326144372792096892477601329560050788540507270643350323540922623768812838108259196176567079601907775012220177855013634617700243158568695595782613158429994895498609846478472911899288934916270337490662530266770655491010497702030941359884700149793050675398807877070203475918458074503234929487127050506598923962668789734434468894649437716320436839496321751776798629259662152088406699583079605572445577680927670146137298092304249370799903292212729601860113190343772421287399409591430084186776240481457300095284459152395320758915322559752935515642817837475136257300083011993342524430843536051600227046970319188710980778393583645738894884897864545557652672823152633565195917603156595268321272593989260122727660622043428814867127758702797028389827674369636792548519994111325778779819588227947944918528217703586639291970443209914849353418633381083317671220838481547988218431135605469566186825129161913417966205448534325656703384212769600427516628546326269553495868366098380944550549245873455772097830380087960407177702871275759516277155122804560151354250683589795537910517895394682695652404298527506417029991004369062511404323527637534558835046067375371108830435200469035703387786891796917993046005596528997743258957246189395932391169259759426267068465958929707002336925548204297240453988771965130651509355657420254959760770992120037534898485938703556174734534905763146988235543622917599990371917782687334363018378938577577742626156399641331467982577709857289285860493677569903899499639049930688104220578029295454192631858805197535815858199098663892456413321679182565758374914970365076277744686231169674078572734292237538026837326139712967052369594856020770609901553667490936264248879718144097755723389654758031500474853517264613170164287929861473663915239675758200752518576500131307233054752205153794844388786082809495574294146831165168782742252201812256714429548940713841777633192318592514717411266641533170529392969154438886064308178666902668860313622225826930040303388269189855873767223121132243089923390781518797892432643417433437316312623054479713120197