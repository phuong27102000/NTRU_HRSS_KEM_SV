`timescale 1ns / 1ps

module Add_in_Rq (v, m1, c);
	input wire [9113:1] v;
	input wire [9113:1] m1;
	output wire [9113:1] c;
	genvar i;
	generate
		for (i=1;i<=701;i=i+1) begin
			carryselectadder entity_0 ( .in1(v[13*i:13*(i-1)+1]), .in2(m1[13*i:13*(i-1)+1]), .cin(1'b0) ,.out(c[13*i:13*(i-1)+1]));
		end
	endgenerate
endmodule
