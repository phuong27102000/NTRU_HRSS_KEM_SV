module Add_in_Rq_test;
	logic [9113:1] v;
	logic [9113:1] m1;
	logic [9113:1] c;
	initial begin
	$monitor("v=%d                m1=%d              c=%d              ",v,m1,c);
	v=9113'd1478487529416704287878515439357116189672197922245827580099170648464021043360570295024381185677859725132159715962919444160031602332326433422338756177122453663543458195597145888663623195797734623057929259245333811391384372678016424552822221788074151479942461363468149136007305662267986090404687836082439124898281076545763023888583914760182570354411989916778496745585078369334770947079273817467766932085848768927569047201455463652914963297803033519868964124496010224818625065721362127361168273907190764913892535236033284011721729262374829119130378885207536053023448308221400590565646052200343352620916790140735192265592176880989229033360340076152329274688598421357141752607864563323313205112161343011489922158467859275550874081173819994162121428753903669002190622878070940925236751714358805147909946270236434537787889071356542940964464324962580121112842532666837867635813915278114971951869803715450953703716826738277018961492041149321307322373647201080486391003375640158504884805160264526431723869840904623476471226332742199758013625413335589872185815163212706443872521982940248258727573754776462305219228866505158481607167790356283648666177634760998174761889823473720902648801241460571311175525582822219162992514410642937939700781361041475902904874234673354780077006933467137869229722538788728367745511877528305004509700382644190290735073193040108078696390790052820192894248383211903140338964992064124075448801770910793059615129708907399907351460739595917186085890285606986986736680057239934152479909543737576755479153911664698159273972112613447689504410047900393725287838125459677527313176820574188469508505183429042114045791324559242023895500804750594423582666459914583338007161868594728841644876221688314150586685567376689762949888207015445333784296007813011528061533038898188623032202451210207461504998581420811680179688692834767640745792054471472174757938531675856393455529130711618581201054526475933914124562257725908875666744383333143181904762898204562990538565214754585134853898708063920280040635821614803747675252787476846387099184552875541633704197738777688883197424684231641015087629523091644051687148583446171940287478719187537478663725357974124953409799637974416265231397179048428155204831269830796179810983521342357035965627378265006518699806361718437126050292393712375228401380998822464022080037813557468590861980401479510631402616612162219111669448103705724847682981407792945198926663363323273533951667316216596510102603186514865610632708931107994319003239678411298904502623844319961690985579125986132297866126267898914424393942352514004119622420905027664531744225364596428646747756265095685732214617992474329657158803539019157912174925386671093355348711332403838609531460527742686231347080713612528857917336534405691672322569058;
	m1=9113'd2360263817128565792877628832464064110429040439711828239654720771964859286615981153602764681509983918753067887052361927967288624714079881584383036351510709769369348906808138572594969892644816963424964494695327124696869940548153814821210795811660016346593518392339514390113621046628513211758098522446996858486877129644648413462108733624636734644303339081258057458047635863222967179095177261733971510349345105104272627294421046220943774109867138621904308495310943370733678189337887693973504636548133356708476206190479023984209931532463550879441563256011619508437777641448345653950466800785146968469988049149106479688863186270316735546361818880949508417606817289898873319817978717004551242246245315704910947209135639596572237639808139347720151919764534933876154285072534424656301118509654755944461803415511550671870149895517835440912756129565716002926426265477462299999607861537236118505526260741889140931119369896986288516322397502266862027464963955979377769490487649867417615760819862951343468995676521803076104460193448533400232900867352042596804626336185674399018537053245044203300244416548589198713010430849600444375481594696827369830076789418283568777659078593372752212323473896016201279599719455283045406908757225542493765120627727472780667758861577498861485738118564143753483169306569645352541612635806251118581714580537199811403591760813239861999263938020427207310050751691395819914792276900201853967302795378884962446148992702098094292163701925121505773906097427159928954751667020497091184082040243402059478580776638303296912131348459537017942882552146406110644329268665866015654535822973554568493583037363719307588443542921973295237988765926329072811434428578748760583858786396136746269945847422580157814510475322036473910499751562707126464123823934891827682184239095156666261118785953675277746326167665271419962978987006046594134528010271571427694463612198476001647662164661645053282444408492218094484246379845926582980038347301995771978566225838837898879469124200414001095989819590948786455414602029547570017329159632726021196300752923266529399240000731245323045477218220776643562911456338272707993095296767110137881817270591129765232776730623480388986697397990289002707015564223477454166656009115470065152522436562217965373816257602900887568714914931052917881447663839465121064189875224237305342024049227063103732091169900710577489546174021053018246968113394623503347060219568645983461408119863971216328886015610738094620181752632747498536647911950773357001971524728763270720046377783127979373241760549885631511554532257751504695165734122064085596332208826339229418656432706373851626778563255469037448564970535067545753657753823465728146658041941096117912060789962656533441548893218208473399365963446071424516133088386805598765057;
	//c=9113'd1480847793198662182596310039167829848087509530108117785343173259227716657924149956472606352051993902686742948426432007899872488444101772221985433507268943894558067747026864814852677680150744030347168393713481511175434191546962653702274938208392101047120133515465257098095282298973476832769892925665602793821896452566244906363587945912833258024294208881751223535448717886201277331806372474015686489616013181249627705566175841056286332604205308611167387743408114087689753546581431212399475797975052046190657586047127520602779928501932715688369293670308218829853207326049609184985510727871023869099453925866889545471076695429758041954038654538365315699399210999218898751244610017542213525956302326846567636292078215412706825376092836439049024049025784269175882012574376245058046595876326155303601650916685259476760005604314277576771011230979666043673634918272577274255442346705854671969010796727531547978897714714315516334488013409071602425365265985131562666192095512598471552452415961717932772066800240491285449379977526128163116886087768382856933846083512927872995753916457744213492468236087009245103062672081463003058991798716148125538549389876227553939020489209432333104874742870874787971508157878781389442212478410428332199248353869551350722814709156343398431819342054379306356341814200289324596049806357978080222997638427749833069739441903683416394292254573822246996932053207961033673358826496345548823536367547439545716883926035201627529058537278271243177977022412682187699605797341110375420949663374251935624323441722591959730945202244922581594347895298365665420089112573244085353039268147740054280659295979943429685187941683988410314551821118612317688569642317924521681898659564396700238171332290713108729768958212046731294269987024794296615874479171694126213914114317080559356146252568724201525669896042553902136839032637256447584491782723351940891690219424885191198746583550948160264088955686360341809638847217502794815521099666344284919827335720256054394105512115060706064405438378478279388157285248763428209978273346791570178243583829420750652091041279377971825411748860294698231031016696671829230604346057019191916339466482364454957524577480666186353232854273700171134756973631900349917118510579837010462776848623429578051744245662653219900096083033524017720440560250492864092900503781195009943014007537101799970222221214702993336357837770805238809914574908456128691331349783358532551644625728220905523536030331711687182112008057883845010014573360314200627300913988932626246910178622746415432030057627887219087519848877696803134156418636548732335494021690341691446702418581826645325260544094283965041929095703272914545770159048964283340646479817793855930301445674252891239330562918478369153834355543031195406650128217922458046870371;
	#20
	v=9113'd9016705096966681476960796913803553018982658760093196142124536481692524306804030018286215530773595474295841874220778381399119480764859964014567930860884046138154280548891675282558559470151603769411778087313175684862654053583287107803451956039155834684917111402319299740706813164781266952221160326612682144777031236366901448163868186112887738962244910811868084104608578437025221755524787311821116888629330849075154563087867633396119504438733310259071968516766718877971454582442001942483307627707873546399105844540190418420485109660597528906406123802712493480016110155960734100867133392336521554313568711185854248040972354913242527273316257253163440832178348641181233300860829468478604370013242932666478609351991112185630739137326484205748652525545508363614447905605155634455630879096229454884531342842523860030091004928615988678085054841148509496092959420671319384532782860613330370441386329598745588179831404536414734812343229851028263789390835243777780494554794797527792994372171356650010544743315105825129202366768214756421412463885199047581656947769835548820818755701231721209234573977652692460389393925614406756757428984197752466828597753160094864654811633985400074923423721007738418252541210150381063856355094012786591548455856085363664939551608336830605910997216715233578062624861613998089105939416645544989815510735602472211611633435434043018842969746014962914982023999462362196621569553624815663989629566915436852912284730363629855024936480119863712984098570361821629173688858017890340577723783692140067231202025904767541894056783051114460710219278133982332513170827844983468810335158874004662415627835099328355946661294716277234196750858068069777817528573945615722384582333644438595541161353693342695224878440152180264558365884784920952629381389219864496163721092805158828051442910628264178962530414488589683921366744899288350909373977052384133744495083703690922632779806368096690012547618707438125522885408068906306045603489997082958383686310577591559916478158392985547451442128607044706770152769049306734405899279044891760031648343559512035680329836497741277755450729265315483509641944030188262696455127101140402029371761098497836962728953388302306585494526348933072017196400335925454862848146815369024126051721320152853168920781026278125279932380305663314122353704168934602346715592584503511252218119334952435885205988395972810064407941170055577215524813930594132464437734273798264257132375848254902504714863036841726647911816671347503055233527387895911837500721997687678380523498139028246322454482787926303097879875455247559354750185469701046257536080650490668632290363789915105146362416007315259740448010483140416832574445626617648209084150555582465215142512060771927803312216965286955617502354812347333228209753309652202788780070;
	m1=9113'd288153303824860447797294346778089477547045093689636546948754091568073861206819203685564133137971465262868918394470732124665836633909449171840629540931584360604742274292590990831099361815856238895964466688896697629749252321337109127538063198390062836973691873753654225437552540446636789814958366754797941402801559764177826710674517622254728628600869008594998726840820579936200986011109735583519489912295702846415521111837630729548971624036659873370913627059889358426579265580583580254024260404294309353326323731131934871345273957286408215933954300935089977437936810743759221778746576486989413390170576914383776063245541727359806801070687831581244761821781247869760835194967815766719463424474879845873233255180705781694238887456985477303276189437950945345625261181405145912205033778361652746641529687693474539294254818787990458448526243654216782517027368543044865605394750730350426573391221746445819162888216716918288352859156745189165127124259423985791845967060545938917991996811704392294631987176146162656399373676163392542851586416471356060103502054851660095231268042126888696469279135649625710039939464108061035248504256226415830339530912406463084567260951238174923275452340693587999567915421666794102289444757435210629622658332398672571898661633917408485369681228307086473527005630723470124151855791894484716989625138806747430292173182677589595589849242317136006558445165630824657467500252481139308562855328655841209029342328436993763851979365052216473405875054816616031334496736288353656673939698777150932949012973283234377394059998692150641773755720963954278097958267488744596384609218831263138333670935587508168997563516774650940896274541678437107146772924315468610403288920719493448898518678203091196747784368932337689148196021879150398797453745760255484724907961328407126008187404162689350873479743708543841437848422669671920175613479769031438883393850931896001600227384476352470050813403090873201018530015768243884878520010329637831794721433783690626296138658689112241305408534503549316852172444670969108296817878946586536499635400283595490067674028399113297735002575842878556824504028729476319070876144327651423951708640595789620044956323455670400591938467041321537416164100513003626037002003237706213264393171836606138897014598011069141071384320343739744668113526770305943170920323859502251438376180032705097801964722087064902627960397789908082694796199353650639449110178123306785696617412297278271739908108837748111853439009646941971381292457028539995283463189906223574779010286861976385002411712405675644159350366485845628498831163912639697834417952299693882750538088208159719460560217181295205199817611392660016936101222043034822697694545102080832631344174166666442515352582387256612742946770358294642638060370956644261888;
	//c=9113'd9016705385084814630746161682077102694312498006650191956014582925818744657401573821539327940216799273422884825326962945096908090997295719066251464966698859933638952407746066997485069285208802168324264100774379306849568695034357999289347459081413461244975744136036311795826247225746140154641494578688142473019686970924555090733848970448871325543038700456718096582171507740062048702499830244206103372899217198653337105512264058065471327110235247924224050733553862825096713519255839644935631064434358223865254342069331542270880742514434221992630591485823828168968823586491203632588363829240178825141654916949965715407394196577225654356077645642736254542724313058993585531793956324423678529916547870224736748910450349080744396199363293444902123055324097717459384238778233468656317931848143493084198435084770050124188797788100528326408456870774693000401424156864714059270004963366437538898658287046892342517110110282973149867934600960673344345171950519407588109431079805338382059234910455567662289111220553127882342762788832238664687119807482403812761377173227396829817333079473799636983377706274710362430193233298694759002607227918027685435065047999128895536972077859417749597725931322076417366614446521844419197796785972442287614220094233088803303671847898571601378360840299405714415385747108308407603000304716999830256731447377046603427712152207205486954034814999642315664364805645994313986266251199173526494939564633291137004685189497601984324964895631391787165345733496186716373471634775914636619139317936249478880201853156720146883640003083557703933148580708842952562507101996232206880135680137417007973059506407713627311302416162203432321061061162657379427716189158891229474414333075184666850054556306859275606630406390582566290568042685518914398043763427694388476836820623707122899508090902849269800138673221403530699658731602030572772024188144476211219036125612863917815095267595805506412445243210428137373711621900541522915774908013184316037957042687662405762940842363289985221738840915214247194921300551848956956934482631857792374557447338782029531560744101562474213903649865822085446546993921546402759548774014488764369302975850829457325721950754372031036241507262036166676613806139442846320402088712782116578323766270858995187099253819316074005814068595022847843555640451288788189260490785446825404246925087492158630210621808516099226266930024061415301792901097618163374598628669504200870522003951685136068604897666649689732779106573569794455064060760783772109887157987846497539772872364295012093207497893953817779936612754854303748029710719049397537389461112051587969920920954175594137678964126777388395046547306823273541760335641975020013979263587423805619790341471157114975694223803603949315078412175414087902516240241710702529124390;
	#20
	v=9113'd10571629790255253433201853975422425973333640877513881973702323624914812374897059179190850573091808548225763945909172207674988554770443571305487282013801641020165920948266158719074712139843409957439269188625922989337293562654566162541382070284254208764631011939949045684229985127506790225193821044463445048569824999984516951891967560225850162587457345156718750691312177578776785493476561787929744075013483647519137495459544831595832164445240501877811624914079465252120282217199576847991563754009967115019175549186160016653427449364088840448525227564572004836288130930502841056288886405037125087395011449362735353578250627969964346707763189289904265117876723627011337333743509045128164799503261651262480373633592758013603001881945363708745940486300556545409919398034323271276104798667051850340439725398214495121821847546840085429359754798612842401474396164344049560192180394764998406530640326250817999741476099330405002167003290933379496470736260840256090572039577344954992210597500273399969516523380054353925499009821059580163225630272167126867978141339599348161670983510097065596728922661655624196069571589012360994391763551117402320566697610575800562799651941506115757650359422207736220201797652381900973843465842375821352487196586256109180073748495903037863372162256697352475696727423428171689287544404295911223961770446781606208153316651691633663375431501095639487459318644381623131175997693328666418826377615673125623527525470730161424931896968170850451959720180870875159598414396169549983739922402160669338393086969298792656308647914004828439036157973675347563914316472651878919202224932727474636458587117066202213065218312346509408179370783218614584417127002582848493413139279697356472358056234690927722391047941003116914886777050713895586067024701836704823860587258782950399543923014817938967685639278114017186517077494270734922902158315195665293910719069240029761905449448433903173177673526242388682030823510425226237529545482344692257713252894222620326044767804785752397375613953080751415036761465439745088806223879444893504114984580335760500323199435435412862737734920080058960060369524093032649909106408350096185262945377707310635562380860529569975809289325346988463071241678688159509361389545474516103533953608926594439216991444044160196862077965741143570163283000747924759435906696699630901187052638620921695472108405684902280260258867717534167024152184185377149695222039185351135926712203913479170599367827529416017731235962533825939086210644270651510328190728345987463217524341415808792276591265817523136281452564699867651219266145523984057845932861599822412624170533375854848799898459324123669226067738925348027271441187602335109438892851145854758185722852560684785758483968501468238360515256548797262112103045516208832856915243;
	m1=9113'd2359975663829034751194690464038648926146261720797916275623434120002745387516974736245380357338286526522408740902739758299964799113895253638143181385311224632634924560175082507965585782095642285906241603138887652833347451052937104143938335179835737691229537754874027325832122398301795960187554388248326020286203612187429648525939811718622373857899697019593407507344465482655374438944190648610773204743923471534647936581878620790798618415813779893175137963099917947587823200820156241095994529804521161298620815922612650132045721899775293328161583634570743085194273016774534106627810001636495923845494390574092068574937272506337458845210915826147358622274012615607915279900371659814850523372781846480329763690192309029752499143712862624716065240612162840280004119205647795505370473551530930264046417006488645015945596617226037735292295817775495562031653703448050676603028658389119119325659542406230476594326199845121099531350441479966369615474229815403820318038797705781292542566470719046864364864045014904080496410561849994548198160466578664325179699217940853493144687581071998707982821795590358131450345387049608253494869204517334966344169920009350705377956652708459383655163076645834771076918595483150354263626474961390664870997031449554308930370836370218181204693354450308480320387533258399045326053739341221958390007677353235360205284303570031405623436835601559916796032226525308855791603689030522584889587778639350445341129218843875772612416757735074251230046284944128726197185466906466592901337191074001805236780152527623856445591476777003604133283081903406784821339865556821260152060239034174913508020063339097358791658542866492054827016906799297329143444292471361817254061760864718863550101228697777813548749767654676929372016976307834515025728452639996709480031049129227955103095575229192675339252486315727873797272261513271497430173308595922617472664655379600569657644833645287897731120940110093614882647729123048115406942387988081411991044080887044019194323516143465757422444836656268265159578904910228196966835391040218953460595786694586315258015992536566063458454529706986265445535744523360254414631447193785691629852998918297340636075714744924773721186911521925851759947284336051536432471261753926270058774246046875615056775739364246034904085952295453154243783614959696211264320388898881849609021553082630986222821773988007034466178566280554446843287748585784922640450172414214471543967336387329717935017205688782419680408611008309437661103118176211735383600511044682418263838996823766023646410187973364440312196302749991682308571100104362135206992465227416828573662147910044043837203648209294760423616002170402822039914514561851400475920996744096343333500232829889846615549650523390058560865314232460206496734313221452214575103;
	//c=9113'd10571629502137115986645700100961119873361740037846531970096733551950494345951774330611831838745264607902505740347718049984662180506607686333183448398769963242882380939664079992359701162541842317430386114269052791474036841912824424581379869130948643524129184615612094011502395528600933573038410768258485511399242996606894702724036101140182591972905800694405306318485987587025001759886047745151072204070303913616799644823282773586162804304731913494667367633958466493103575746260640767054198244561749130121548894156199076496688733816058512037713420158834815845006209926336787750314061462072606004836558112544588484627043534726516319167442234144122011856083270023398210800163350276245098500906266286868732520009062281711615776548750994866035076318193314867074635511075262668873803154536746983661320523965476054805070256701595709479727305511804327360878902646306650556519871532164206801334178218001241222889578243710839628900392985632989051925875146820461402060966721772252609396010445114772354802781442823775752139826418832722306497305116433103156678865494402021978099749870164304002027145141081956275853098097456121369165414624700895931533090748507172774966558546428147507111132783545438000323041064937649632128782628728315826920311519289048059862415264496502828370727271116050016556139076145790051574592302326673300354294194595629416957644799848925346689965282689143286117195226095292574683334229154721260105490974573481170378585706305510874575279372123416016459886971204248107121217661448344264379431930519293963094948529346654315973199644915931533216564246626586429310149680344940838020145081431745281959820224644018901289053253242316341442551545927838094362517205670565615528141793105850977280050067908229678388624469136816924923640021809194008124423071375213924137433586090492447930191308394783287902579494728120073794434948086870493112079297379200017381094585434962946796722372928939367286612071676276711036484619115177046266870617132613127200760132190836936627426931241377733821172530912822985500549558787010764816923953611826448372756695412894738213723872654811239133857772242034195302369202545345580442555240976582147616486037113379602171494300883014220270626284820722143485760699667702478689679018025072844395010118396709712642121952518609896631936369163927328452866256082826508500449299735954468429012947774745644083592080484782080607381748480576039681977604271062865403766877884692987679821304389624066683607717007796895951835839372211045179527708566277740337238944234771293300856718335056882324527605221328496583352071398380165332754981986622764952570360091076420260816103338502301670061083853765821551920723628114036495817550762334957253747301225147290336121048350301159291664413710938082167703886667029866410686755774402239264652586;
	#20
	v=9113'd13551964423202356714105278302060484102970972282232158670204233075434854480706443671994636839432782652274870242857492362267572997450734293256639736733432048088994184592825759756918002368656507473497781379925250425497456908038981470315502710197565048487054097171408965627287820488493706421501784792379516311852778896210189147132495467478074237629022440316792646674962924763813539576097546787968890373655996184439561592745809479936958720204816134001108569151651744143232373892754984994356123401842700067323407244134122247889284087490606205967806808248012763403918971381085857020955198726601055154928691786231385809470584090605111110445267784090526466786395808358748032306213778395326484174012072351765700032392763571933642528303978840657083857353599783899201979620111965178798844961957371829961854749247437326761268264580422815103237722800911397250097315125633874211775994597259704393569873572415914180161252958579973726206913514319420164304129040980142821900909091859618783805304534566714386782596798981980484851938328710033207614992639074820096525106692623122750730240362293708871393940264051156240288114174672783758164023934776335648573914840420110471170495613954823418656872710272172658473578488844003411028534644088074315422279243740609194376695111510569956005712744816607740833753227458317664800327632653710390263913760193782201748056126767438111420915227197104400055555954981393931894932273110494792395777430272424097749390931029409998598401682984795607563049181332358835078354868157958053732034518951030501912156912027020560504297530837292591413276597643200746811195963524927560170215968312702365097663115047849725731038868349612362092122504699112553237288298571516110919733013173443166531752462423818636929834166614594989800742272395708198755660897755462079602910035130248707798322002627112952373505728315933175275301385913301574697455374436246195787275629636069686564373941854254452723324052848368577734809392141620186473903339961967569702284927301202275040134006184375114089052592992965243861662936051155872546363251611671544769842038032775967788198706873632013234884485194889549495157733984826518081465771323582110364584203317846549690495179401115354980123415458400064674555162995230247824396680164670943549095058861096249763572394172895613709286663826737154552187393333495232082951498178647718091592189458119989368909879721929998416638604953606018284958588427938847997565350018687308825102258955240460205600297849233409703268300965984833584067010455959319513249930323145181442438560208278745736495955398789586396711467243525123356992944900207808435374050661000942410013217729224517728749788233875075307698415963228716879079458119575223921811258108174757347466232040259118928678048421729477901610313402835622479176551383554913289019543;
	m1=9113'd2359975699003997549027090047921953566231270431171285518441395043102455852700266284391904298893855237836129381016716133772575179455589680754757331496343991568882689091588947353159591612667378591717459208271966123784362941682478869541068886781512552369012291051484514666666402616320169105127714665315013907108481622973225317715248571546910277543879056036880384963914436776914588468970838877110352492551675724673091287085468449581388188403804897884332156321947731610412290529865627506793790206951827983882810503526251470707946439600267696171277051765586845102248954388417612106656521642267754094173152764436080051382589521907085273285717813620529080949861748593039019735591663479417283088466439480505236423390476223337929887863184890511212952605970749838535369102828345791048995909931914392299338937614451959308006095429778279302369701661911754250084658411098874060631806611746732868097017890527090753982890709401943014956563336972049555924916653429125572017864466473037860419053462875548260429405208072037455126605497923851494339060492773376287421706291454034651476090622433462289947508767397230592297256590968388429081762741102015858198902480963021316115367674805598901606203640019843570347933372898187234443405592630731612410321091511809470178785138642978266660847749221296895898425513071845888940245763130841627289037222017903196030594858172500248146850977037018224979697961642067990755041843370235413689383944514235383220185215996496606919899482881977402099258880231185044503326146930160595211387698007602444855655688905623023490808923108234281394624948238842184276844526805870690655280377765280092087710961958042566219556050513407100845878184110341887245270309459887059468793377424250986876660010351513313284289840368781458982780661678120833082302088184179088490427508551058476740046825201407134312952401516826390723278335124670402271171851937069127495578445802886955979014832391157540925974918564346707061378871273043109054915540698918091985519300365534254626583952918127050140476565061816515979447472177592990028600025737120513486083553638518045634959879544136714588524168534848014973415502453268796124934191041817899029862572858636086255015275103825780905614182392571712755137154511234803637791866829465786826899723801773679447853221933550620740656227655157686526639377151148834200939164042903142143332248117034696087642196407237661889749045007898556160580434218745810689917270234007169398138398600086267277317570742490251014615874490704907753705401827726057044877254544836635172132706001966816042271993910842468143518904865644700215065298113887386307153909944943122574228583996228928998990442963619770328767873757894179402945737377225089260930491832361942885589784788090832568444135871712731725179277209461690295823061965740875710464;
	//c=9113'd13551964135119389937576167720994351580033210286591434455686953881424113950071295318206208259528333619484337906640322231334312879218733470740217903940049143403988688857895523791727960276030127830393019718243544605897543641321071889172405774339226938912993949563586954253775483855704825364062242445015791509788829993204949215121049295917188641569206917768971803755904311097004717404877520048648952899693606290444544335203244593251826580315440721652606202001951230306592984837185651388998046680564173629894536776661130531872313567953559957092729363779780876519772465871276610411385539540530762020248640126160478704283049157610559506954128201741529096401236086596332309851038119216257773121497025846707406734191203994132004858372285939060676279630219326033826633061783293339538052354841630446564122907303041156678268928782291957936677112264288260082705521845855794102023472698053221305417278594270657168889385754168533986386083607776018621175567458806962399117185950165295565642848508294932828388000476497465136893829976873358172279348342044335851130081445048490695902308782881098055078287166708266870708466998892960493088502048499129515284253472164764947420526068626879690419048265966942318287267727032762169381257952417374407938667474056533595434865898710484538276285733049610696525133128985775968791552726783491132583253117462384155230150563507769338823562310947724197886855532585324855406535634710212098202717657353565659304293928028484115957610601438467535563925573636862664866089932207123005195989583920708473712632723583786111613375392460957175092506979144495126198271148147217278033872000218376110636988068042032722282882121971284165421660540994588427992316608672113065296998301115976223204889274183608260753394132722447042398430278972976514406711456548780906638420018093546822922846618550877164004699399201296904027347217296886265747532879340984019590533684611981244036719041079997836679195099171004767147643979966605085846905126965082395696751546959199736622832076945807811054362254729484037966989077443612187995918419864640184526103747593234401796784267153369260111104028392018049396377212422787298336113185808959724181533666843663264704743093238875038518630889307230710593523613193679480902910197428490632090441106451752665817553829528376659818782897313127963846273455273981109864068837567544077562539160964295114121089725031743332015025863916958988033551556073946355243811339483568445510069451652240990360868970215376044097184702013399740796989788935841971017810402324619732824922795360078270855941042436887170227059998478584269444486496145745697669406191169599969216715506817942400433073915782762111341021367646417880106694127317932430428455115980867531965972159924526574005488574406107648178634639015631461911971996328441286824468631;
	#20
	v=9113'd6079418929106854942101211075895337144656737721594258488224651608735830693378563565441886636281139974375827455930240286442658833834382185592019601991926335515129742990722993512379462993534049880861750706403259091324496773909859800661565831015391253511610916907405306537488510189425611876449111206208321493896750083998316592805547681655926642474727740488122175339038989650544895554683385777426409398462190107364356823666805329500116088490628150527246717050390751632242872308175607957585490047910415562946537205636868403483896789043312798417146090514610728990383786933716155955030889353036999566417272899826644536106281931027389175340309449211938010159259643997339516627098040931635911525405441013124252416475463586721838802813376457536041192137821549489086324799160016313133399235745786876720508730285177946247485851894836568229450274637005803260626484506197391767369617950403402227714707346596934094193827957827364740718795797223132418639151619940898216834204401543885269621183950693594633316484690989272234632418746512369502375006861185614292069598580500284736726407240679859089348904161941704003819704263020690168901447651697069000097601936472740439318995367365746803711285009342054079323555689304170151730502744425744391920718021777575574408120287787855999596076231223551765125194584070444635514603045670318681751600666715763551278957790230370745891108372900547675145843532690887071670766363203396188281522380313061082690225282581640848582100607806757837063398294646430061787371688241789355975506286496415857791465001579261246393698648374081834506640996242070616735890025365015821862478152548962458942090647974229722846306565831599117201843183329366192303371379929503507664002319344357188979550969331230160383427913705904033965339222780962626985916783258496166657746433957266153330720161162601108974627119196688420528560728250807138510156567915777378678211644899172791699198323853427879197570232754155612488966440353160837842670149750410809702029145628932736367029741789205811531946064638909678317982915320925248386191243880064927357848090810482205393030220833386104234094465773123461079865702716179484286380178841373213740194873854015606214858410883052430081761466130545778226859030726417871462351363482508250727687030565192143316263914234018220490480606016163303113727041111481765635993638257002498813202494792866572473136985683578787500923029802816359531569338581785481887935617727457279604021727514423112622369991562909081215176224441199706070085489738589043847526443970646275674847021739097848863093527493030684981392199229890601456435103562579795357970936752292245454468586911165140599596685414987941845070717326565480985844763750298756174392201683090333562168746796380492550424392944411912350251726880067106969627260590117966589556817;
	m1=9113'd4720527528775169851789494162971246119510518529748696805310790136935262101649096946517033360686938256772203019354577095363490543098073159732653250684725711125576312952912403331729738461161472575228984583512628105324861345085409597673152058934809287970480197605959935331826045905337249977157745635502980057363173207335726537090221670463754017717512991496025332212809059193096204025520021068477279470224195207019809975295562556611182393863689396849377963240676373895265101813322258009847283473195565048348934553251558583091442309155674051929016942411647273643317423474089555608724236223861996169618244729185204712515228665769716530127712982751335277808994821952288773642245843395845775152407916044893480294572920161118596088304169993716389162327319273719730473536633580436592015022285511006254985027291871438873298414551618681825260505278187068531823311871624882982782877916519712492835534805582694814383956107257460098204277427450723454729662669223039025537920775488389811829913905493065353463479904153207796729120615276369313933056334436638354306273269932883975961901558403906884715892564213334956745444839975921476949748675801568179624921743716984799691379328723290467909561208900648322401596408095708523360850331183092714420433815715224336461090728101723568561073935687898223095237647874095640220803883939270743821328266646646546496386271041733617238692336752926106235201025300527884546519726698767670887772377570636155039636627077253619503168713818068892738200064659340511438566998027761572541066376020246429174549342506760914578820664255394247649288092540116207591850164312452841463948996832649663962527956883446913644238403869460563041856497501408169047453159508115964544362178451840375973247489867888037871880488288938950279223053705948668420203067619462191253519718692285210943315701510993183238402565507659198790031819123097141413697001561421214930892823467956190388873275059708020723342778613214335147657484592183831065107957085115487364235514283148069095995832244976975985459419290090183146438121356148530737598694971338726407839328877618073749229794361774852173156775147271163617415856274280313105713312959836606980257334799302240341847107507558053291795535027497763096330481705071941639350075444213056272255889131948998395115406880754352503542058384028676143025246149988585491378095834355149781540935779891755577048980659317335038171274019305101619749100220763985316316012748003910820560608245329973900121175540297626780156647883259690367360855880348659467331721305813316635878753730152204063175563345819508981809731341027308266206172550855062032862564440092161959694750995154531728792718076180569258347547053956641974517582201055809062666642476605984587308820617477014498284626258290926535231523043985137679109323697278286831616;
	//c=9113'd6081778904735521890794753135651436093521299759157250092920321736458178619616574715769316019861058577797506979526771404460462487970262364366539270131551823524731556752680638865398435290133819266859126096799441964621552791360198428271645811287367202625726077220667041384170381167614764371139516484132398958863189383939027532139678924916724922686793832110276071384623559187162038845611498545367718436979951473357824404982170212821640977529057716628676203796737125151193701891814080215323907083101521320114918569991379873318442478359637614455216926777472367790970761737395888686036306429026481567520375774990182390006183307106699191538198449470285870758204243446185400005471328633594965025154205528227859232743264198846140452722949999137374058844496378311853474656548457874848279576477298723236036715778066053416413618412077184492517529363525159306301302050503215801052330724196916277097729642354868360399108933047480749214964377548425905957679371491073144838996933027530727533080939827411424452812345204283062157089742370529178524841708717292878799299285759902376273640014192041697309499807092122152751796285794098385945455385678735716848380467053828650900871874760572540613246097724147211099754574484373331571333129268670285163686408854835829351000901675594550626466008116241848264358667858720383797921795072097038795790797067869461124380430077084855467884251773795880647993514444813422331183325521402916023984474987023437819001353826304418649143488383056443810098220261571943883371300499258628754231504100974458599138481980828530291007137750127786887076109431279582294503195617478318946171295215999348342078549314654273859155226670838287608615785425487944620319342723173678390865115206724617497029733656330874949523972804561206375887546994127066085757156098591550801991764190345987608192663568534318456774888409098761361622801211808282933279303205689392732950132133991706609490769313582776814925862625135035462468037793040543445652028092183199989349243581189616200826374531917261232103480279115406578285452983833499486973861333619200434971308005419327513883378029125275089587947472402601004034839972852588157269610305569033837441282731206850748185019915048902830225604634181906863074947235285095970817723492334917809953160944551327923317946545314810952787781244454827455045981498913473778744488433949094441502074379911094645853195170063818170346247731250476305079834592911479645794184307760162269445622624963956221333630127018714531683632492572539460652753191051059910350726731190459597387828587179718643626374046727664968644501695962675631039262627273780567162349718458507159263327990009293609904059762498337388576195240867143789613252106446793380132048482132405753650566895220349021353235562457045894016437941181896569701130204700923336693841;
	end
	Add_in_Rq entity_0 (.v(v),.m1(m1),.c(c));
endmodule

