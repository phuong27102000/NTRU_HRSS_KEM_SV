module vector_mul #(parameter NUMS_OF_A = 700*13,parameter NUMS_PARALLEL = NUMS_OF_A/100, parameter NUMS_PARALLEL_2=(NUMS_OF_A+13-13*3)/2)
(
input logic clk,
input logic en,
input logic [NUMS_OF_A:1] v,
output logic [NUMS_OF_A+13:1] b_out
);
//11=1111111111111
//01=0000000000001
//00=0000000000000
logic [NUMS_OF_A+13:1]b_temp,b_temp_3,b_out_2;
logic [NUMS_PARALLEL:1]b_temp_2;
logic [NUMS_OF_A:1] a_S3_out_mod,a_S3_out_mod_1,a_S3_out_mod_2,a_S3_out;
logic [NUMS_OF_A+13:1] a,m,n,a_temp,a_S3_temp,a_temp_2;
logic [NUMS_PARALLEL:1]a1,a2,a3,a4,a6,a7,a9;
logic [13:1]t1,t2,t3,t4,t5,t6,t7,t8,t9;
logic [NUMS_PARALLEL_2+13*3:1] k1,k2,k3;
logic [NUMS_OF_A:1] z1,z2,z3;
assign z1=9100'd2359975699003997548963130587883005460920122192262842660440347650815524605726626959954220389796157611024673610638994781033202834896508335518424008842866055679802473270756462288129033653311516062666649491449942201904195649033552101503599021565654767605657949809025902774084083313848733206875778162950121072934262986237902546156442416052128997203628049572845513012203053118841435494329207026114609879984225950778165073799947308385051192485608328203639298349561753984904653922611197255548117232435639819101740127044302513772603311248422041878137373248377023118842253276447831702176723742191122582701990355946422966093538011485503878963279265863596892835636197820872846401958935899367161090364927030045609105090118878564960962974111195397390107059854729289822174167753935841945116395997207940376995680955448172461901332127472184790828524538590484674163200282203380642498860800398807512831054648576006700346964015483360691267181870580836203568946758399489168213376494899403280039682178547845388272244220530453078685890445393863714558675656017594048363397245253514692554919074973872472240192512496781120332370268013683805331969295331656779770451420782379654436644277991736324598306245515452029248960809707895038562344558900459125975346580872614874507456863474538130800574184999355335099398268892064290739918841782886502279421465484484232713048451106001574036094738699047665922789173547338217056668888098021790111206630719751124597989564058323040193723887894435895849649427507870999749029021967144392171293538230143713987201419736693778917724592917694403970053141717198090211985467296028748833850750269629304905810249796490477803360544842792697365085665985676531179928172988412412281495026688639205543193241341748727743908819661181161232561684363073910419763888328261859921713632138095972122768564905365890577653763988965830777939640736741855519137168868950763060180363392374277700343627964562610064453699052137652581766911210803013486791358358064755490338442086455713296356795885510860336203909377579308415784387153489423492265186985434184077003011261148911080353169542567962520867003750458060458997828161899969939050555314427086772959936727333604108714315529196591026437097188536910080410665087846967699690952121951999430345964639749532286077226476982029832925761846990649829656796219509017395807456137671451586570419840077468063840926310118521895538910959016283318394404979373749961680205200514307897827078412397520082334941720368374225971507429897918101958268789591741468939357056804883726182432096222071176357834993567291158581163232152486820938885619828710186395058981997920686550779575642295045191473688344901606893357828914904171931186961662215152403476218600805892137888100859328073345263168757632416842763560575405341880681942160938893313;
assign z2=9100'd19332920926240747921105965775937580735857640999017207074327327955480777570112528055944973433210123149514126218354645246223997623472196284566929480440758728128941861034036939064353043687927939585365192633957926517999170756882858815517483184665843856225549924835540195525296810507048822430726374710887391829477482383260897658113576272299040745092120982100750442595967411149549039569544863957930884136830778988774728284569168350290339368842103424644213132079609888644338924934030927917450176368112761398081455120746926192825166325747073367065701361650704573389555738840660637304231720896029676197494704995913096938238263390089247776467183745954585746109531732548590357724847602887615783652269482230133629788898253853204160208683918912695419757034329942342223250782240242417214393516009127447568348618387031428807895712788252137806467273020133250450744936711810094223350667676867031145111999681134646889242329214839690782860753883798210179636811844808615266003980246215911670085076406663949420726224654585471620594814528666531549664670974096130444192950233116792361409897062185963292591657062373630937762777235568097733279492467356932339879538039049254129144989925308303971109324763262583023607486953127076155902726626512561159990039190508461051965086625583416367518303723514718905134270618763790669741415151885406226673020645248894834385292911460364894503688099422598479239488909699794674128231531298994504591004718856201212706730508765782345266986089631218858800328110144479229944045747954846860667236665181337304983154030482995436893999865181752557322675336947286755016584948089067510446905346208803265788397566332849994165129583352157776814781775754662143425971593121074481410007258633332371809839033071605577678101050664396072817145318302301474158705773185121156478678074475282203629720083704757375612139634597608085732881536915389280412771687374444650988997536910330082921215000285696901648004702635111649949834536638898286483794807669266476976852517572245203323754871894104967874182425621129694542105699561385357248636411784676835958808668251331879570253164892716748970942494723752431280110208302284553740702149135786694844087801670316884858587672815178473688572700168494367378724168399642359395868279783030779333394142328828168487544639299436788391327841050547403404548474630217870506454680679804531397184879329914618378984868332490931368254758576261392944286965591029759686084241002613210298999426354360484514487842573257721659158588865723745091242137924335546113551213009345607484886483732251207076723384267303249171096889197793172037131350997636793846948323180526966264223986283661681010208552454921433963670387334470894976460283589936866528489277182777801868393579322239615576844395878462524758775919088233720560686546470182411414020096;
assign z3=9100'd2360551864937550607184277103139129634152494890547905313812890334183479200222139897698644652700728488487911664944195088226886062616761969927611869329941406350639210245318871406815579909402100269715341909959201161991698713766188503682856328853337091692078303425058508920064840398846188745770224705950747145394323246680305997452842004170414576503737153317723039876861562734925209503514898815964494240146364735727842819956666045569787982064981090018302945895772840729947892282389797637595557937784478282339158397152580559862850763571960907872671401937605742365707823071748912637370101893381119961270008951020888378698722229827161279695238786462345245840954540785818988432006188797827709061813475068224096631859926184781824856284025417712313834348459637025624255718518950448832334127729931787431096851345280360165313351074330024045752888007925452287974348518332443845511525313281295789285080651225085527645239905570210467197809853602762902555808879525995610727800627929178436311715546580517293115146107741341855946515420903072724658647383940455272507904546598640442302517503446955327591587256834736154975812441682055211503990078506158221825528864419573232860201685628498188737427017864695592501197586468459492759722405297974502928447008459799509404847254154188093233272512873036414856967888833744902456151573911610267042262837916733411803998927261822224564977799290844827165317205005995159210912592177186864848468979594023234550197707559929997966628096839277427451661958096370968187764183288668928287832192480948116713870619219359571516946811810807110451042347452401538009205813296511389938857195480557622528987695177882794196481887343271263801643386254446076202729800974019891540875859598127509594409070304889835548563785108154986216154797140247335741451743411601986566780776438149211353548190537887932555078388686272029752125849080651450957578069530266203985794505514512067218748115939121605391938356031626846662198779689073795882177178348761746216861300126318596899554351251761753809567845570043778991667692822127776251195790979423862582962995646558579645992121414532739213375241980131852314206781169285577611085998628045728787705670047824550288978542654265803052882720059206815457677705129538786633084605821634889610220433672164875971794216485772938973475261102096144834535650976087509488174072456802070942949918397682399225735857558495305860517812414137763318353897742469763928214821703117714355344757902714284806497824721784218068649059490139051416587561410238200438266597106205052597889610362565246452260225630586157114869856143117316071445816017147139972192788966855793720651154021529122023475735110312494483020310042761601118773204130473710536490408904766459080178565470561242650453864480420044320435037786389047274955044539011442941951;
integer dem,dem1,dem2,dem3;
genvar i;
generate 
	for (i=1;i<=NUMS_OF_A/2-1;i=i+13) begin
		mul_in_S3 entity_0 (a1[i+12:i],a2[i+12:i],a3[i+12:i]);
		mul_in_S3 entity_1 (a4[i+12:i],a2[i+12:i],a6[i+12:i]);
		mul_in_S3 entity_2 (a7[i+12:i],a2[i+12:i],a9[i+12:i]);
	end
endgenerate
genvar j;
generate
	for (j=40;j<40+NUMS_PARALLEL_2-1;j=j+13) begin
		sub_in_S3_3 entity_0 (k1[j-27:j-39],k2[j+12:j],k2[j-1:j-13],k2[j-14:j-26],k1[j+12:j]);
	end
endgenerate
N_13_bit_adder N_13_bit_adder (a3,t1);
adder_13_bit adder_13_bit (t1,t2,1'b0,a[13:1]);
N_13_bit_adder N_13_bit_adder_1 (a6,t4);
adder_13_bit adder_13_bit_1 (t4,t5,1'b0,a[26:14]);
N_13_bit_adder N_13_bit_adder_2 (a9,t7);
adder_13_bit adder_13_bit_2 (t7,t8,1'b0,a[39:27]);
//S3
genvar o;
generate 
	for(o=1;o<NUMS_PARALLEL;o=o+13) begin
		adder_13_bit entity_0 ( a_S3_temp[o+12:o], ~a[NUMS_OF_A+13:NUMS_OF_A+1],1'b1,a_S3_out[o+12:o]);
		mod3 entity_1 ({a_S3_out[o+12],1'b0,a_S3_out[o+11:o]},a_S3_out_mod[o+12:o]);
	end
endgenerate
//
//
genvar p;
generate
	for(p=14;p<=NUMS_PARALLEL+13;p=p+13) begin
		adder_13_bit entity_2 (b_temp[p-1:p-13],~b_temp[p+12:p],1'b1,b_temp_2[p-1:p-13]);
	end	
endgenerate
//
always @(posedge clk) begin

if (en==1) begin
	dem=0;
	dem1=0;
	dem2=0;
	dem3=0;
	a_temp=0;
	a[NUMS_OF_A+13:40]=0;
	a_S3_out_mod_1=0;
	a_S3_out_mod_2=0;
	//k1=0;k2=0;k3=0;
end
else begin
	if (dem==NUMS_OF_A/NUMS_PARALLEL) begin
		dem=NUMS_OF_A;
		a_temp_2=a;
	end
	else if (dem==NUMS_OF_A) begin 
		if (dem1==3) begin
			a[NUMS_OF_A+13:40]=m[NUMS_OF_A+13:40];
			dem1=dem1+1;
		end
		else if (dem1==4) begin
			if (dem2==NUMS_OF_A/NUMS_PARALLEL+1) begin 
				if (dem3==NUMS_OF_A/NUMS_PARALLEL+1) begin
				b_out[NUMS_OF_A+13:NUMS_OF_A+1]=a_S3_out_mod_1[NUMS_OF_A:NUMS_OF_A-12];
				b_out[13:1]=~a_S3_out_mod_1[13:1]+1;
				end
				else begin
					b_temp=a_S3_out_mod_1>>(dem3*NUMS_PARALLEL);
					b_out=b_out_2;
					if (dem3 !=0) begin
					b_out[NUMS_OF_A+13:NUMS_OF_A-NUMS_PARALLEL+14]=b_temp_2;
					b_out_2=b_out>>NUMS_PARALLEL;
					end
					dem3=dem3+1;
				end 
			end
				
			else begin
				a_S3_temp=a>>(dem2*NUMS_PARALLEL);
				
				a_S3_out_mod_1=a_S3_out_mod_2;
				if (dem2 != 0) begin
				a_S3_out_mod_1[NUMS_OF_A:NUMS_OF_A-NUMS_PARALLEL+1]=a_S3_out_mod[NUMS_PARALLEL:1];
				a_S3_out_mod_2=a_S3_out_mod_1>>NUMS_PARALLEL; 
				end
				dem2=dem2+1;
			end
		end
		else begin
			m=n;
			if (dem1!=0) begin
			a_temp_2=k1;
			a_temp_2[40+NUMS_PARALLEL_2-1:40]=k1[40+NUMS_PARALLEL_2-1:40];
			k1[39:1]=a_temp_2>>(NUMS_PARALLEL_2);
			end
			else k1[39:1]=a_temp_2[39:1];
			k2=v>>(NUMS_PARALLEL_2*dem1);
			if (dem1!=0) begin
			m[NUMS_OF_A+13:NUMS_OF_A+13-NUMS_PARALLEL_2+1]=k1[40+NUMS_PARALLEL_2-1:40];
			n=m>>NUMS_PARALLEL_2;	
			end
			dem1=dem1+1;
	end
	
	end
 
	else begin
		if (dem!=0) a_temp=a;
		else ;
		a2=v>>(NUMS_PARALLEL*dem);
		a1=z1>>(NUMS_PARALLEL*dem);
		a4=z2>>(NUMS_PARALLEL*dem);
		a7=z3>>(NUMS_PARALLEL*dem);
		t2=a_temp[13:1];
		t5=a_temp[26:14];
		t8=a_temp[39:27];
		dem=dem+1;
		
		
	end
		
end
end

endmodule
module sub_in_S3_3(
input logic [12:0]a,b,c,d,
output logic [12:0]e);
logic [12:0] t,t1;
adder_13_bit entity_0(a,~b,1'b1,t);
adder_13_bit entity_1(t,~c,1'b1,t1);
adder_13_bit entity_2(t1,~d,1'b1,e);
endmodule
module mul_in_S3(
input logic [12:0] a,
input logic [12:0] b,
output logic [12:0]c);
always_comb begin
	if ((a==13'd0)||(b==13'd0))
		c=13'd0;
	else if ((a==13'd1)&&(b==13'd1) || (a==13'd8191)&&(b==13'd8191))
		c=13'd1;
	else  
		c=13'd8191;
end
endmodule
module N_13_bit_adder #(parameter N=7*13)
(
input logic [N:1] A,
output logic [13:1] S		
);
logic [N+13:1] B;
assign B[13:1]=13'd0;
assign S=B[N+13:N+1];

genvar i;
generate
	for (i=1; i<=N-1; i=i+13) begin
		adder_13_bit entity_0 ( B[i+12:i], A[i+12:i],1'b0,B[i+25:i+13]);
	end
endgenerate
endmodule

module adder_13_bit(
    input logic [12:0] A,
    input logic [12:0] B,
    input logic C,
    output logic [12:0] S
    );

    assign S=A+B+C;

endmodule
