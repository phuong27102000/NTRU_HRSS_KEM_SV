`timescale 1ns / 1ps

module sub_ter (x, y, z);
    input [1:0] x,y;
    output [1:0] z;

    assign z[0] = (x[1] ^ y[1]) | (x[0] ^ y[0]);
    assign z[1] = ( x[1] & (~y[0]) ) | ( (~x[0]) & (~y[1]) & y[0] )
    | ((~x[1]) & x[0] & y[1]);

endmodule // sub_ter

module sub_2i2_o13 (x, y, z);
    input [1:0] x;
    input [1:0] y;
    output [12:0] z;

    assign z[0] = x[0] ^ y[0];
    assign z[1] = ( x[1] & (~y[1]) ) | ( (~x[0]) & (~y[1]) & y[0] )
    | ((~x[1]) & x[0] & y[1]);
    assign z[2] = ( x[1] & (~y[1]) ) | ( (~x[0]) & (~y[1]) & y[0] );
    assign z[12:3] = {10{z[2]}};

endmodule // sub_2i2_o3

module add_ter (x, y, z);
    input [1:0] x,y;
    output [1:0] z;

    assign z[1] = ( x[1] ^ y[0] ) & ( x[0] ^ y[1] );
    assign z[0] = (x[0] ^ y[0]) | (x[1]&y[1]) | ( (~(x[1]|y[1])) & y[0] );

endmodule // add_ter

module mul_ter (x, y, z);
    input [1:0] x,y;
    output [1:0] z;

    assign z[1] = (x[1] & (~y[1]) & y[0]) | ((~x[1]) & y[1] & x[0]);
    assign z[0] = x[0] & y[0];

endmodule // mul_ter

module inverse_phi1 (clk, rst, z);
    input clk, rst;
    output reg [1402:1] z;

    always @ ( posedge clk ) begin
        if (rst) begin
            #0.2 z <= 1402'b0001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001110001;
        end else begin
            #0.2 z <= {z[1398:1],z[1402:1399]};
        end
    end
endmodule // inverse_phi1
